module main (SW, KEY);  // keyboard selection keys are missing + sounddevices output
	output KEY[3:0];    // KEY0 is our record button. KEY0 again is stop recording. KEY3 is total reset (of saved recordings).
	output SW[2:0];    // SW2,1,0 are our registers for saved recordings
	
	// simply call the music player module:
	
	
	// simply call the recording saver module:
	
	
	// simply call the recording player module:
	
endmodule